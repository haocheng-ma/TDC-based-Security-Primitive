`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
module TDC(
            input wire	clk_delay,
			input wire	clk_sample,
			output [63:0] data,
			input wire	ena
    );


endmodule
